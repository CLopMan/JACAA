package Constants is
    constant WORD_SIZE: positive := 32;
    constant REG_ADDR_SIZE: positive := 5;
end package Constants;
