package Constants is
    -- Sizeo of CPU registers
    constant WORD_SIZE: positive := 32;
    -- Size of register IDs
    constant REG_ADDR_SIZE: positive := 5;
    -- Size of a microaddress
    constant MICROADDRESS_SIZE: positive := 12;
    -- Size of the operation code in a instruction
    constant OPCODE_SIZE: positive := 7;
end package Constants;
