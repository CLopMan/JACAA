use library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity StateRegister is 
    generic(constant SIZE: integer := 32);

    port(
        
    );

end StateRegister;