library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_std.all;
use Work.Constants;
use Work.Types;


entity CPU is
end CPU;


architecture Rtl of CPU is
    signal internal_bus: Types.word := (others => '0');
begin
    

end Rtl;
